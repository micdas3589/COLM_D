LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY KEY_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		KEY_RD1	:IN STD_LOGIC;
		KEY_RD3	:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DATA_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		KEY1		:OUT STD_LOGIC_VECTOR(127 downto 0);
		KEY3		:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE ARCH_KEY_REG OF KEY_REG IS
	TYPE MEMORY_BLOCK IS ARRAY (0 to 15) OF STD_LOGIC_VECTOR(0 to 127);
	CONSTANT SBOX	:MEMORY_BLOCK :=
	(
		 X"637c777bf26b6fc53001672bfed7ab76"
		,X"ca82c97dfa5947f0add4a2af9ca472c0"
		,X"b7fd9326363ff7cc34a5e5f171d83115"
		,X"04c723c31896059a071280e2eb27b275"
		,X"09832c1a1b6e5aa0523bd6b329e32f84"
		,X"53d100ed20fcb15b6acbbe394a4c58cf"
		,X"d0efaafb434d338545f9027f503c9fa8"
		,X"51a3408f929d38f5bcb6da2110fff3d2"
		,X"cd0c13ec5f974417c4a77e3d645d1973"
		,X"60814fdc222a908846eeb814de5e0bdb"
		,X"e0323a0a4906245cc2d3ac629195e479"
		,X"e7c8376d8dd54ea96c56f4ea657aae08"
		,X"ba78252e1ca6b4c6e8dd741f4bbd8b8a"
		,X"703eb5664803f60e613557b986c11d9e"
		,X"e1f8981169d98e949b1e87e9ce5528df"
		,X"8ca1890dbfe6426841992d0fb054bb16"
	);
	SIGNAL GEN_KEYS	:MEMORY_BLOCK;
	SIGNAL KEYS_POS1	:STD_LOGIC_VECTOR(3 downto 0) := (OTHERS => '0');
	SIGNAL KEYS_POS3	:STD_LOGIC_VECTOR(3 downto 0) := (OTHERS => '0');
	SIGNAL COUNTER 	:STD_LOGIC_VECTOR(3 downto 0) := (OTHERS => '0');
	SIGNAL PREV_KEY	:STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL CUR_KEY		:STD_LOGIC_VECTOR(31 downto 0) := (OTHERS => '0');
	SIGNAL RND_CONST	:STD_LOGIC_VECTOR(7 downto 0) := (OTHERS => '0');
	SIGNAL RUN_GEN		:STD_LOGIC := '0';
BEGIN
	PROCESS(CLK, INIT, GEN_KEYS, KEYS_POS1, KEYS_POS3)
	BEGIN
		IF INIT = '1' THEN
			COUNTER		<= X"F";
			RND_CONST	<= X"01";
			RUN_GEN		<= '0';
			KEYS_POS1	<= X"0";
			KEYS_POS3	<= X"0";
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				IF ADDR_WR = X"0" THEN
					PREV_KEY(127 downto 96)	<= DATA_WR;
				END IF;
				IF ADDR_WR = X"1" THEN
					PREV_KEY(95 downto 64)	<= DATA_WR;
				END IF;
				IF ADDR_WR = X"2" THEN
					PREV_KEY(63 downto 32)	<= DATA_WR;
				END IF;
				IF ADDR_WR = X"3" THEN
					PREV_KEY(31 downto 0)	<= DATA_WR;
					GEN_KEYS(CONV_INTEGER(KEYS_POS1)) <= PREV_KEY(127 downto 32) & DATA_WR;
					KEYS_POS1	<= KEYS_POS1 + 1;
					KEYS_POS3	<= KEYS_POS3 + 1;
					RUN_GEN	<= '1';
				END IF;
			END IF;
			
			IF KEYS_POS1 = X"B" THEN
				RUN_GEN		<= '0';
				KEYS_POS1	<= X"A";
				KEYS_POS3	<= X"A";
			END IF;
			
			IF RUN_GEN = '1' THEN
				COUNTER	<= COUNTER + 1;
			ELSE
				COUNTER	<= X"F";
			END IF;
		
			IF COUNTER = X"0" THEN
				CUR_KEY(7  downto  0) <= SBOX(CONV_INTEGER(PREV_KEY(31 downto 28)))(CONV_INTEGER(PREV_KEY(27 downto 24) & "000") to CONV_INTEGER(PREV_KEY(27 downto 24) & "000")+7);
				CUR_KEY(31 downto 24) <= SBOX(CONV_INTEGER(PREV_KEY(23 downto 20)))(CONV_INTEGER(PREV_KEY(19 downto 16) & "000") to CONV_INTEGER(PREV_KEY(19 downto 16) & "000")+7);
				CUR_KEY(23 downto 16) <= SBOX(CONV_INTEGER(PREV_KEY(15 downto 12)))(CONV_INTEGER(PREV_KEY(11 downto  8) & "000") to CONV_INTEGER(PREV_KEY(11 downto  8) & "000")+7);
				CUR_KEY(15 downto  8) <= SBOX(CONV_INTEGER(PREV_KEY(7  downto  4)))(CONV_INTEGER(PREV_KEY(3  downto  0) & "000") to CONV_INTEGER(PREV_KEY(3  downto  0) & "000")+7);
			END IF;
			IF COUNTER = X"1" THEN
				CUR_KEY(31 downto 24)	<= CUR_KEY(31 downto 24) XOR RND_CONST;
				
				IF RND_CONST(7) = '1' THEN
					RND_CONST	<= (RND_CONST(6 downto 0) & '0') XOR X"1B";
				ELSE
					RND_CONST	<= RND_CONST(6 downto 0) & '0';
				END IF;
			END IF;
			IF COUNTER = X"2" THEN
				PREV_KEY(127 downto 96)	<= CUR_KEY XOR PREV_KEY(127 downto 96);
				PREV_KEY(95  downto 64)	<= CUR_KEY XOR PREV_KEY(127 downto 96) XOR PREV_KEY(95 downto 64);
				PREV_KEY(63  downto 32)	<= CUR_KEY XOR PREV_KEY(127 downto 96) XOR PREV_KEY(95 downto 64) XOR PREV_KEY(63 downto 32);
				PREV_KEY(31  downto  0)	<= CUR_KEY XOR PREV_KEY(127 downto 96) XOR PREV_KEY(95 downto 64) XOR PREV_KEY(63 downto 32) XOR PREV_KEY(31 downto 0);
			END IF;
			IF COUNTER = X"3" THEN
				GEN_KEYS(CONV_INTEGER(KEYS_POS1)) <= PREV_KEY;
				KEYS_POS1	<= KEYS_POS1 + 1;
				KEYS_POS3	<= KEYS_POS3 + 1;
				COUNTER		<= (OTHERS => '0');
			END IF;
			
			IF KEY_RD1 = '1' THEN
				KEYS_POS1	<= KEYS_POS1 - 1;
				IF KEYS_POS1 = X"0" THEN
					KEYS_POS1	<= X"A";
				END IF;
			END IF;
			IF KEY_RD3 = '1' THEN
				KEYS_POS3	<= KEYS_POS3 - 1;
				IF KEYS_POS3 = X"0" THEN
					KEYS_POS3	<= X"A";
				END IF;
			END IF;
			
			KEY1	<= GEN_KEYS(CONV_INTEGER(KEYS_POS1));
			KEY3	<= GEN_KEYS(CONV_INTEGER(KEYS_POS3));
		END IF;
	END PROCESS;
END ARCHITECTURE;