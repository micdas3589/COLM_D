LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY OR32 IS
	PORT
	(
		DIN1	:IN STD_LOGIC_VECTOR(31 downto 0);
		DIN2	:IN STD_LOGIC_VECTOR(31 downto 0);
		DOUT	:OUT STD_LOGIC_VECTOR(31 downto 0)
	);
END ENTITY;

ARCHITECTURE OR32_ARCH OF OR32 IS
BEGIN
	DOUT	<= DIN1 OR DIN2;
END ARCHITECTURE;