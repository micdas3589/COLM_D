LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY KEY_REG_TB IS END ENTITY;

ARCHITECTURE ARCH_KEY_REG_TB OF KEY_REG_TB IS
	COMPONENT KEY_REG IS PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		KEY_RD1	:IN STD_LOGIC;
		KEY_RD3	:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DATA_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		KEY1		:OUT STD_LOGIC_VECTOR(127 downto 0);
		KEY3		:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
	END COMPONENT;

	SIGNAL CLK		: STD_LOGIC := '0';
	SIGNAL INIT		: STD_LOGIC := '0';
	SIGNAL WR			: STD_LOGIC := '0';
	SIGNAL KEY_RD1	: STD_LOGIC := '0';
	SIGNAL KEY_RD3	: STD_LOGIC := '0';
	SIGNAL ADDR_WR	: STD_LOGIC_VECTOR(31 downto 0) := (OTHERS => '0');
	SIGNAL DATA_WR	: STD_LOGIC_VECTOR(31 downto 0) := (OTHERS => '0');
	SIGNAL KEY1		: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL KEY3		: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	
	SIGNAL CLKp :time := 40 ns;
BEGIN
	tb: KEY_REG PORT MAP (CLK, INIT, WR, KEY_RD1, KEY_RD3, ADDR_WR, DATA_WR, KEY1, KEY3);

	PROCESS
	BEGIN
		CLK <= '0'; wait for CLKp / 2;
		CLK <= '1'; wait for CLKp / 2;
	END PROCESS;

	PROCESS
	BEGIN
		INIT <= '1'; WR <= '0';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00000000"; wait for CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00010203"; wait for CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000001"; DATA_WR <= X"04050607"; wait for CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000002"; DATA_WR <= X"08090A0B"; wait for CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000003"; DATA_WR <= X"0C0D0E0F"; wait for CLKp;
		INIT <= '0'; WR <= '0';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00000000"; wait for 45*CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '1'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00000000"; wait for 12*CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00000000"; wait for CLKp;
		INIT <= '0'; WR <= '1';	KEY_RD1 <= '0'; KEY_RD3	<= '0'; ADDR_WR <= X"00000000"; DATA_WR <= X"00000000"; wait for CLKp;
		
		wait;
	END PROCESS;
END ARCHITECTURE;