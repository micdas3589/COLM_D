-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.0 Build 145 04/22/2015 Patches 0.01we SJ Web Edition"
-- CREATED		"Sun Nov 05 17:17:26 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY COLM_D IS 
	PORT
	(
		INIT :  IN  STD_LOGIC;
		WR :  IN  STD_LOGIC;
		RD :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		ADDR_WR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DIN :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DOUT :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COLM_D;

ARCHITECTURE bdf_type OF COLM_D IS 

COMPONENT control
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 DRL_CTX : IN STD_LOGIC;
		 DRL_PTX : IN STD_LOGIC;
		 DRL_TAG : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 TAG_CTR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TAG_INTVL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TAG_LEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 WR_PTX : OUT STD_LOGIC;
		 WR_CTX : OUT STD_LOGIC;
		 WR_TAG : OUT STD_LOGIC;
		 RD_PTX : OUT STD_LOGIC;
		 RD_CTX : OUT STD_LOGIC;
		 RD_TAG : OUT STD_LOGIC;
		 DBL_L : OUT STD_LOGIC;
		 DBL_L2 : OUT STD_LOGIC;
		 WR_RO : OUT STD_LOGIC;
		 INIT_DK1 : OUT STD_LOGIC;
		 INIT_DK3 : OUT STD_LOGIC;
		 KEY_RD1 : OUT STD_LOGIC;
		 KEY_RD3 : OUT STD_LOGIC;
		 RUN_DK1 : OUT STD_LOGIC;
		 RUN_DK3 : OUT STD_LOGIC;
		 TAG_VER : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT ctx_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 CTX_CTR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 TAG_CTR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tag_ver_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 VERIFY : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 STATE : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 TAG : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 TAG_VER : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or32
	PORT(DIN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT key_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 KEY_RD1 : IN STD_LOGIC;
		 KEY_RD3 : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 KEY1 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 KEY3 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT l_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 DBL_L : IN STD_LOGIC;
		 DBL_L2 : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 CTX_CTR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 LA : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LC2 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mem_out
	PORT(CLK : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mem_out_32
	PORT(CLK : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT params_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 TAG_INTVL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TAG_LEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ptx_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ro_inv
	PORT(INPUT1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 INPUT2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 OUTPUT1 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 OUTPUT2 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ro_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR_RO : IN STD_LOGIC;
		 IV_WR : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 IV_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RO_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 RO : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT round
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 RUN : IN STD_LOGIC;
		 ROUND_KEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_OUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tag_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT xor128
	PORT(DIN1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	CTX_CTR :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	DBL_L :  STD_LOGIC;
SIGNAL	DBL_L2 :  STD_LOGIC;
SIGNAL	DRL_CTX :  STD_LOGIC;
SIGNAL	DRL_PTX :  STD_LOGIC;
SIGNAL	DRL_TAG :  STD_LOGIC;
SIGNAL	INIT_DK1 :  STD_LOGIC;
SIGNAL	INIT_DK3 :  STD_LOGIC;
SIGNAL	KEY1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	KEY3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	KEY_RD1 :  STD_LOGIC;
SIGNAL	KEY_RD3 :  STD_LOGIC;
SIGNAL	LA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LC2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	PTX :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	PTX_OUT :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	RD_CTX :  STD_LOGIC;
SIGNAL	RD_PTX :  STD_LOGIC;
SIGNAL	RD_TAG :  STD_LOGIC;
SIGNAL	RO_IN :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	RUN_DK1 :  STD_LOGIC;
SIGNAL	RUN_DK3 :  STD_LOGIC;
SIGNAL	STATE_IN3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUTA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUTB :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	TAG_CTR :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	TAG_INTVL :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	TAG_LEN :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	TAG_VALID :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	TAG_VER :  STD_LOGIC;
SIGNAL	WR_CTX :  STD_LOGIC;
SIGNAL	WR_PTX :  STD_LOGIC;
SIGNAL	WR_RO :  STD_LOGIC;
SIGNAL	WR_TAG :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(127 DOWNTO 0);


BEGIN 



b2v_CONTROL : control
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 RD => RD,
		 DRL_CTX => DRL_CTX,
		 DRL_PTX => DRL_PTX,
		 DRL_TAG => DRL_TAG,
		 ADDR_WR => ADDR_WR,
		 TAG_CTR => TAG_CTR,
		 TAG_INTVL => TAG_INTVL,
		 TAG_LEN => TAG_LEN,
		 WR_PTX => WR_PTX,
		 WR_CTX => WR_CTX,
		 WR_TAG => WR_TAG,
		 RD_PTX => RD_PTX,
		 RD_CTX => RD_CTX,
		 RD_TAG => RD_TAG,
		 DBL_L => DBL_L,
		 DBL_L2 => DBL_L2,
		 WR_RO => WR_RO,
		 INIT_DK1 => INIT_DK1,
		 INIT_DK3 => INIT_DK3,
		 KEY_RD1 => KEY_RD1,
		 KEY_RD3 => KEY_RD3,
		 RUN_DK1 => RUN_DK1,
		 RUN_DK3 => RUN_DK3,
		 TAG_VER => TAG_VER);


b2v_CTX_MEMORY : ctx_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_CTX,
		 LOAD => RD_CTX,
		 DIN => DIN,
		 DRL => DRL_CTX,
		 CTX_CTR => CTX_CTR,
		 DOUT => SYNTHESIZED_WIRE_0,
		 TAG_CTR => TAG_CTR);


b2v_inst : tag_ver_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 RD => RD,
		 VERIFY => TAG_VER,
		 ADDR_WR => ADDR_WR,
		 STATE => RO_IN,
		 TAG => STATE_OUTB,
		 TAG_VER => TAG_VALID);


b2v_inst1 : or32
PORT MAP(DIN1 => TAG_VALID,
		 DIN2 => PTX_OUT,
		 DOUT => DOUT);


b2v_KEY_REG : key_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 KEY_RD1 => KEY_RD1,
		 KEY_RD3 => KEY_RD3,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 KEY1 => KEY1,
		 KEY3 => KEY3);


b2v_L_REG : l_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 DBL_L => DBL_L,
		 DBL_L2 => DBL_L2,
		 ADDR_WR => ADDR_WR,
		 CTX_CTR => CTX_CTR,
		 DATA_WR => DIN,
		 LA => LA,
		 LC2 => LC2);


b2v_MEM_OUT_CTX : mem_out
PORT MAP(CLK => CLK,
		 LOAD => RD_CTX,
		 DIN => SYNTHESIZED_WIRE_0,
		 DOUT => SYNTHESIZED_WIRE_6);


b2v_MEM_OUT_PTX : mem_out_32
PORT MAP(CLK => CLK,
		 LOAD => RD_PTX,
		 DIN => SYNTHESIZED_WIRE_1,
		 DOUT => PTX_OUT);


b2v_MEM_OUT_TAG : mem_out
PORT MAP(CLK => CLK,
		 LOAD => RD_TAG,
		 DIN => SYNTHESIZED_WIRE_2,
		 DOUT => SYNTHESIZED_WIRE_8);


b2v_PARAMS_REG : params_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 TAG_INTVL => TAG_INTVL,
		 TAG_LEN => TAG_LEN);


b2v_PTX_MEMORY : ptx_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_PTX,
		 LOAD => RD_PTX,
		 DIN => PTX,
		 DRL => DRL_PTX,
		 DOUT => SYNTHESIZED_WIRE_1);


b2v_RO_INV : ro_inv
PORT MAP(INPUT1 => STATE_OUTA,
		 INPUT2 => SYNTHESIZED_WIRE_3,
		 OUTPUT1 => STATE_IN3,
		 OUTPUT2 => RO_IN);


b2v_RO_REG : ro_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR_RO => WR_RO,
		 IV_WR => WR,
		 ADDR_WR => ADDR_WR,
		 IV_IN => DIN,
		 RO_IN => RO_IN,
		 RO => SYNTHESIZED_WIRE_3);


b2v_ROUND_CTX : round
PORT MAP(CLK => CLK,
		 INIT => INIT_DK1,
		 RUN => RUN_DK1,
		 ROUND_KEY => KEY1,
		 STATE_IN => SYNTHESIZED_WIRE_4,
		 STATE_OUT => STATE_OUTA);


b2v_ROUND_PTX : round
PORT MAP(CLK => CLK,
		 INIT => INIT_DK3,
		 RUN => RUN_DK3,
		 ROUND_KEY => KEY3,
		 STATE_IN => STATE_IN3,
		 STATE_OUT => SYNTHESIZED_WIRE_7);


b2v_ROUND_TAG : round
PORT MAP(CLK => CLK,
		 INIT => INIT_DK1,
		 RUN => RUN_DK1,
		 ROUND_KEY => KEY1,
		 STATE_IN => SYNTHESIZED_WIRE_5,
		 STATE_OUT => STATE_OUTB);


b2v_TAG_MEMORY : tag_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_TAG,
		 LOAD => RD_TAG,
		 DIN => DIN,
		 DRL => DRL_TAG,
		 DOUT => SYNTHESIZED_WIRE_2);


b2v_XOR128_CTX : xor128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_6,
		 DIN2 => LC2,
		 DOUT => SYNTHESIZED_WIRE_4);


b2v_XOR128_PTX : xor128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_7,
		 DIN2 => LA,
		 DOUT => PTX);


b2v_XOR128_TAG : xor128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_8,
		 DIN2 => LC2,
		 DOUT => SYNTHESIZED_WIRE_5);


END bdf_type;