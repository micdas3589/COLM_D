LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TAG_VER_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		RD			:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		VERIFY	:IN STD_LOGIC;
		TAG		:IN STD_LOGIC_VECTOR(127 downto 0);
		STATE		:IN STD_LOGIC_VECTOR(127 downto 0);
		TAG_VER	:OUT STD_LOGIC_VECTOR(31 downto 0)
	);
END ENTITY;

ARCHITECTURE TAG_VER_REG_ARCH OF TAG_VER_REG IS
	SIGNAL TAG_VALID	:STD_LOGIC;
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			TAG_VALID	<= '1';
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF VERIFY = '1' AND STATE /= TAG THEN
				TAG_VALID	<= '0';
			END IF;
		END IF;
	END PROCESS;
	
	TAG_VER	<= X"00000001"
					WHEN TAG_VALID = '1' AND RD = '1' AND ADDR_WR = X"00000010"
					ELSE (OTHERS => '0');
END ARCHITECTURE;
